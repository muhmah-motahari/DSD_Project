library ieee;
use ieee.std_logic_1164.all;

entity CoolHeatSystems is
	port(chs_conf	:	in	std_logic_vector(7 downto 0);
			chs_power	:	out	std_logic_vector(3 downto 0);
			chs_mode	:	out	std_logic);
end entity;

architecture struct of CoolHeatSystems is

begin 

end architecture;
