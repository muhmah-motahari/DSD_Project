library ieee;
use ieee.std_logic_1164.all;

entity DanceLight is
	port(clk,	load,	din	:	in	std_logic;
			p	:	in	std_logic_vector(7 downto 0);
			q	:	out	std_logic_vector(7 downto 0));
end entity;

architecture struct of DanceLight is

begin

end architecture;
